
class packet_type2 extends uvm_sequence_item;

   `uvm_object_utils(packet_type2)


endclass
