`ifndef WB_SVTB_SLAVE_MON
 `define WB_SVTB_SLAVE_MON

class wb_svtb_slave_mon;


   task run();
   endtask

endclass


`endif
