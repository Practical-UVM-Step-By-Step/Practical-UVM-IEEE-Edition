`ifndef WB_ENV__SV
 `define WB_ENV__SV

 `include "mstr_slv_src.incl"
 `include "wb_env_cfg.sv"
 `include "wb_env_cov.sv"

`endif // WB_ENV__SV
