`include "wb_env_top.sv"
`include "wb_master_if.sv"
`include "wb_slave_if.sv"
`include "wb_svtb_config.sv"
`include "wb_svtb_transaction.sv"
`include "wb_svtb_gen.sv"
`include "wb_svtb_master_mon.sv"
`include "wb_svtb_slave_mon.sv"
`include "wb_svtb_master.sv"
`include "wb_svtb_slave.sv"
`include "wb_svtb_scoreboard.sv"
`include "wb_svtb_env.sv"
`include "test1.sv"
