`ifndef WB_TEST_PKG
 `define WB_TEST_PKG

package wb_eth_test;
   import uvm_pkg::*;
 `include "eth_blk_env.sv"
 `include "eth_blk_env_test.sv"
 `include "eth_blk_base_test.sv"
 `include "eth_blk_env_test.sv"  
 `include "eth_transmit.sv"  
 `include "eth_transmit_barrier.sv"  
 `include "eth_transmit_virt_sequence_test.sv"  
 `include "eth_transmit_event_sync.sv"
 `include "eth_transmit_event_callback.sv"
 `include "eth_transmit_event_heartbeat.sv"
 `include "eth_transmit_event_sync.sv"
 `include "eth_transmit.sv"
 `include "eth_transmit_virt_sequence_test.sv"
endpackage
`endif
