value of v in inst00.u1.v is           7
value of v in inst01.u1.v is           7
value of v in inst02.u1.v is           7
value of v in inst03.u1.v is           7
value of v in inst04.u1.v is           7
value of v in tom05.u1.v is           7
value of v in tom06.u1.v is           7
value of v in tom07.u1.v is           7
value of v in tom08.u1.v is           7
value of v in tom09.u1.v is           7
value of v in tomm10.u1.v is           7
value of v in tomm11.u1.v is           7
value of v in tommm12.u1.v is           7
value of v in tommm13.u1.v is           7
value of v in tommmm14.u1.v is           7
value of v in tomm15.u1.v is           7
value of v in tommommomm16.u1.v is           7
value of v in tommommommomm17.u1.v is           7
value of v in TOMMMM18.u1.v is           7
value of v in TOMMMM19.u1.v is           7
value of v in tom20.u1.v is           7
value of v in tom21.u1.v is           7
value of v in tom22.u1.v is           7
value of v in tom23.u1.v is           7
value of v in tom24.u1.v is           7
value of v in a.u1.v is           7
value of v in aa.u1.v is           7
value of v in aaa.u1.v is           7
value of v in aaaaa.u1.v is           7
value of v in b.u1.v is           7
value of v in ab.u1.v is           7
value of v in aaaaab.u1.v is           7
value of v in abc.u1.v is           7
value of v in abbc.u1.v is           7
value of v in abbbc.u1.v is           7
value of v in aaaaabbbb.u1.v is           7
value of v in aaabbbccc.u1.v is           7
value of v in abd.u1.v is           7
value of v in abcdef.u1.v is           7
value of v in abcdefabc.u1.v is           7
value of v in cab.u1.v is           7
value of v in caab.u1.v is           7
value of v in cb.u1.v is           7
value of v in def.u1.v is           7
