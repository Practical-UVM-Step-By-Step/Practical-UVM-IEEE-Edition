`include "class_A.sv"
`include "class_P.sv"
